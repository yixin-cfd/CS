`ifndef ISNEG_V
`define ISNEG_V


module IsNeg(input[15:0] in, output out);
  // your code here
  assign out = in[15];
endmodule

`endif 